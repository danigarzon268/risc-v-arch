module test();
  logic [31:0] A = 4'b00000000000000000000000000000001;
  logic [31:0] B = 4'b00000000000000000000000000000100;
  logic [31:0] Adder_Result;
  
  
  ADDER internADDER(A, B, Adder_Result);
  
  

  initial
    begin
      $dumpfile("outTB_ADDER.vcd");
      $dumpvars(1);
      
      #50 A = 4'b00000000000000000000000000000001;
      #50 A = 4'b00000000000000000000000000000010;
      #50 A = 4'b00000000000000000000000000000011;
      #50 A = 4'b00000000000000000000000000000100;
      #50 A = 4'b00000000000000000000000000000101;
      #50 A = 4'b00000000000000000000000000000111;
      
      
      #50 $finish;
      
    end
  
  
endmodule